
`ifndef REGISTERS_IF_VH
`define REGISTERS_IF_VH

